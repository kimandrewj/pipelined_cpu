module inputMux (A, B, );